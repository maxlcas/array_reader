module reader

pub struct Reader {
	bytes []u8
mut:
	offset int
}
