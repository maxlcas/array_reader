module reader

pub fn (mut reader Reader) read_ascii() {
	// not implemented
}
